typedef enum { 
    Add,
    Sub,
    And,
    Or,
    Xor,
    Not,
    Sll,
    Sra,
    Srl,
    Eq,
    Neq
} alu_ops;
