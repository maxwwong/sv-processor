typedef enum { 
    Add,
    Sub,
    And,
    Or,
    Xor,
    Sll,
    Sra,
    Srl,
    Eq,
    Neq,
    Slt,
    Sltu
} alu_ops;
