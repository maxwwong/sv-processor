module decode (
    input logic[31:0] 
    output
);

    always_comb begin : decoder

endmodule